package count_pkg;

//	parameter int no_of_transactions=1;

	`include "count_trans.sv"
	`include "count_gen.sv"
	`include "count_drv.sv"
	`include "count_wr_mon.sv"
	`include "count_rd_mon.sv"
	`include "count_rm.sv"
	`include "count_sb.sv"
	`include "count_env.sv"
	`include "count_test.sv"
endpackage
